library verilog;
use verilog.vl_types.all;
entity ContadorCarrosPeaje_vlg_vec_tst is
end ContadorCarrosPeaje_vlg_vec_tst;
